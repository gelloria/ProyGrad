`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/09/2016 08:26:15 PM
// Design Name: 
// Module Name: Deco_Sum
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Deco_Sum (Input, Output);
	input [7:0]Input;
	output reg[3:0]Output;
	
	
	always @ (Input)
		case(Input)
			8'd0: Output=4'd0;
                  8'd1: Output=4'd1;
                  8'd2: Output=4'd1;
                  8'd3: Output=4'd2;
                  8'd4: Output=4'd1;
                  8'd5: Output=4'd2;
                  8'd6: Output=4'd2;
                  8'd7: Output=4'd3;
                  8'd8: Output=4'd1;
                  8'd9: Output=4'd2;
                  8'd10: Output=4'd2;
                  8'd11: Output=4'd3;
                  8'd12: Output=4'd2;
                  8'd13: Output=4'd3;
                  8'd14: Output=4'd3;
                  8'd15: Output=4'd4;
                  8'd16: Output=4'd1;
                  8'd17: Output=4'd2;
                  8'd18: Output=4'd2;
                  8'd19: Output=4'd3;
                  8'd20: Output=4'd2;
                  8'd21: Output=4'd3;
                  8'd22: Output=4'd3;
                  8'd23: Output=4'd4;
                  8'd24: Output=4'd2;
                  8'd25: Output=4'd3;
                  8'd26: Output=4'd3;
                  8'd27: Output=4'd4;
                  8'd28: Output=4'd3;
                  8'd29: Output=4'd4;
                  8'd30: Output=4'd4;
                  8'd31: Output=4'd5;
                  8'd32: Output=4'd1;
                  8'd33: Output=4'd2;
                  8'd34: Output=4'd2;
                  8'd35: Output=4'd3;
                  8'd36: Output=4'd2;
                  8'd37: Output=4'd3;
                  8'd38: Output=4'd3;
                  8'd39: Output=4'd4;
                  8'd40: Output=4'd2;
                  8'd41: Output=4'd3;
                  8'd42: Output=4'd3;
                  8'd43: Output=4'd4;
                  8'd44: Output=4'd3;
                  8'd45: Output=4'd4;
                  8'd46: Output=4'd4;
                  8'd47: Output=4'd5;
                  8'd48: Output=4'd2;
                  8'd49: Output=4'd3;
                  8'd50: Output=4'd3;
                  8'd51: Output=4'd4;
                  8'd52: Output=4'd3;
                  8'd53: Output=4'd4;
                  8'd54: Output=4'd4;
                  8'd55: Output=4'd5;
                  8'd56: Output=4'd3;
                  8'd57: Output=4'd4;
                  8'd58: Output=4'd4;
                  8'd59: Output=4'd5;
                  8'd60: Output=4'd4;
                  8'd61: Output=4'd5;
                  8'd62: Output=4'd5;
                  8'd63: Output=4'd6;
                  8'd64: Output=4'd1;
                  8'd65: Output=4'd2;
                  8'd66: Output=4'd2;
                  8'd67: Output=4'd3;
                  8'd68: Output=4'd2;
                  8'd69: Output=4'd3;
                  8'd70: Output=4'd3;
                  8'd71: Output=4'd4;
                  8'd72: Output=4'd2;
                  8'd73: Output=4'd3;
                  8'd74: Output=4'd3;
                  8'd75: Output=4'd4;
                  8'd76: Output=4'd3;
                  8'd77: Output=4'd4;
                  8'd78: Output=4'd4;
                  8'd79: Output=4'd5;
                  8'd80: Output=4'd2;
                  8'd81: Output=4'd3;
                  8'd82: Output=4'd3;
                  8'd83: Output=4'd4;
                  8'd84: Output=4'd3;
                  8'd85: Output=4'd4;
                  8'd86: Output=4'd4;
                  8'd87: Output=4'd5;
                  8'd88: Output=4'd3;
                  8'd89: Output=4'd4;
                  8'd90: Output=4'd4;
                  8'd91: Output=4'd5;
                  8'd92: Output=4'd4;
                  8'd93: Output=4'd5;
                  8'd94: Output=4'd5;
                  8'd95: Output=4'd6;
                  8'd96: Output=4'd2;
                  8'd97: Output=4'd3;
                  8'd98: Output=4'd3;
                  8'd99: Output=4'd4;
                  8'd100: Output=4'd3;
                  8'd101: Output=4'd4;
                  8'd102: Output=4'd4;
                  8'd103: Output=4'd5;
                  8'd104: Output=4'd3;
                  8'd105: Output=4'd4;
                  8'd106: Output=4'd4;
                  8'd107: Output=4'd5;
                  8'd108: Output=4'd4;
                  8'd109: Output=4'd5;
                  8'd110: Output=4'd5;
                  8'd111: Output=4'd6;
                  8'd112: Output=4'd3;
                  8'd113: Output=4'd4;
                  8'd114: Output=4'd4;
                  8'd115: Output=4'd5;
                  8'd116: Output=4'd4;
                  8'd117: Output=4'd5;
                  8'd118: Output=4'd5;
                  8'd119: Output=4'd6;
                  8'd120: Output=4'd4;
                  8'd121: Output=4'd5;
                  8'd122: Output=4'd5;
                  8'd123: Output=4'd6;
                  8'd124: Output=4'd5;
                  8'd125: Output=4'd6;
                  8'd126: Output=4'd6;
                  8'd127: Output=4'd7;
                  8'd128: Output=4'd1;
                  8'd129: Output=4'd2;
                  8'd130: Output=4'd2;
                  8'd131: Output=4'd3;
                  8'd132: Output=4'd2;
                  8'd133: Output=4'd3;
                  8'd134: Output=4'd3;
                  8'd135: Output=4'd4;
                  8'd136: Output=4'd2;
                  8'd137: Output=4'd3;
                  8'd138: Output=4'd3;
                  8'd139: Output=4'd4;
                  8'd140: Output=4'd3;
                  8'd141: Output=4'd4;
                  8'd142: Output=4'd4;
                  8'd143: Output=4'd5;
                  8'd144: Output=4'd2;
                  8'd145: Output=4'd3;
                  8'd146: Output=4'd3;
                  8'd147: Output=4'd4;
                  8'd148: Output=4'd3;
                  8'd149: Output=4'd4;
                  8'd150: Output=4'd4;
                  8'd151: Output=4'd5;
                  8'd152: Output=4'd3;
                  8'd153: Output=4'd4;
                  8'd154: Output=4'd4;
                  8'd155: Output=4'd5;
                  8'd156: Output=4'd4;
                  8'd157: Output=4'd5;
                  8'd158: Output=4'd5;
                  8'd159: Output=4'd6;
                  8'd160: Output=4'd2;
                  8'd161: Output=4'd3;
                  8'd162: Output=4'd3;
                  8'd163: Output=4'd4;
                  8'd164: Output=4'd3;
                  8'd165: Output=4'd4;
                  8'd166: Output=4'd4;
                  8'd167: Output=4'd5;
                  8'd168: Output=4'd3;
                  8'd169: Output=4'd4;
                  8'd170: Output=4'd4;
                  8'd171: Output=4'd5;
                  8'd172: Output=4'd4;
                  8'd173: Output=4'd5;
                  8'd174: Output=4'd5;
                  8'd175: Output=4'd6;
                  8'd176: Output=4'd3;
                  8'd177: Output=4'd4;
                  8'd178: Output=4'd4;
                  8'd179: Output=4'd5;
                  8'd180: Output=4'd4;
                  8'd181: Output=4'd5;
                  8'd182: Output=4'd5;
                  8'd183: Output=4'd6;
                  8'd184: Output=4'd4;
                  8'd185: Output=4'd5;
                  8'd186: Output=4'd5;
                  8'd187: Output=4'd6;
                  8'd188: Output=4'd5;
                  8'd189: Output=4'd6;
                  8'd190: Output=4'd6;
                  8'd191: Output=4'd7;
                  8'd192: Output=4'd2;
                  8'd193: Output=4'd3;
                  8'd194: Output=4'd3;
                  8'd195: Output=4'd4;
                  8'd196: Output=4'd3;
                  8'd197: Output=4'd4;
                  8'd198: Output=4'd4;
                  8'd199: Output=4'd5;
                  8'd200: Output=4'd3;
                  8'd201: Output=4'd4;
                  8'd202: Output=4'd4;
                  8'd203: Output=4'd5;
                  8'd204: Output=4'd4;
                  8'd205: Output=4'd5;
                  8'd206: Output=4'd5;
                  8'd207: Output=4'd6;
                  8'd208: Output=4'd3;
                  8'd209: Output=4'd4;
                  8'd210: Output=4'd4;
                  8'd211: Output=4'd5;
                  8'd212: Output=4'd4;
                  8'd213: Output=4'd5;
                  8'd214: Output=4'd5;
                  8'd215: Output=4'd6;
                  8'd216: Output=4'd4;
                  8'd217: Output=4'd5;
                  8'd218: Output=4'd5;
                  8'd219: Output=4'd6;
                  8'd220: Output=4'd5;
                  8'd221: Output=4'd6;
                  8'd222: Output=4'd6;
                  8'd223: Output=4'd7;
                  8'd224: Output=4'd3;
                  8'd225: Output=4'd4;
                  8'd226: Output=4'd4;
                  8'd227: Output=4'd5;
                  8'd228: Output=4'd4;
                  8'd229: Output=4'd5;
                  8'd230: Output=4'd5;
                  8'd231: Output=4'd6;
                  8'd232: Output=4'd4;
                  8'd233: Output=4'd5;
                  8'd234: Output=4'd5;
                  8'd235: Output=4'd6;
                  8'd236: Output=4'd5;
                  8'd237: Output=4'd6;
                  8'd238: Output=4'd6;
                  8'd239: Output=4'd7;
                  8'd240: Output=4'd4;
                  8'd241: Output=4'd5;
                  8'd242: Output=4'd5;
                  8'd243: Output=4'd6;
                  8'd244: Output=4'd5;
                  8'd245: Output=4'd6;
                  8'd246: Output=4'd6;
                  8'd247: Output=4'd7;
                  8'd248: Output=4'd5;
                  8'd249: Output=4'd6;
                  8'd250: Output=4'd6;
                  8'd251: Output=4'd7;
                  8'd252: Output=4'd6;
                  8'd253: Output=4'd7;
                  8'd254: Output=4'd7;
                  8'd255: Output=4'd8;
                  default: Output=4'd0;
			
		endcase

endmodule
